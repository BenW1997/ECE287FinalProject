module randomGen(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36);

input in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15;
output out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36;

assign out1 = in1;
assign out2 = in2;
assign out3 = in3;
assign out4 = in4;
assign out5 = in5;
assign out6 = in6;
assign out7 = in7;
assign out8 = in8;
assign out9 = in9;
assign out10 = in10;
assign out11 = in11;
assign out12 = in12;
assign out13 = in13;
assign out14 = in14;
assign out15 = in15;
assign out16 = 1'b0;
assign out17 = in8;
assign out18 = in3;
assign out19 = in13;
assign out20 = in6;
assign out21 = in11;
assign out22 = in9;
assign out23 = in1;
assign out24 = in4;
assign out25 = in5;
assign out26 = in2;
assign out27 = in7;
assign out28 = in10;
assign out29 = in12;
assign out30 = in14;
assign out31 = 1'b0;
assign out32 = in15;
assign out33 = 1'b0;
assign out34 = 1'b0;
assign out35 = 1'b0;
assign out36 = 1'b0;

endmodule

